   // GPIO
   input [`GPIO_INPUT_W-1:0] gpio_input,
   output [`GPIO_OUTPUT_W-1:0] gpio_output,
   output [`GPIO_OUTPUT_W-1:0] gpio_output_enable,
   //output [1:0] SENSOR_OUTPUT,
   input [1:0] SENSOR_IN,
   output GPIO_SENSOR_OUTPUT_I,
   output GPIO_SENSOR_OUTPUT_O,			     
			  

